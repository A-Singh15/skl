configuration cfg_sram of async is
	for Behavioral
	end for;
end cfg_sram;

